/*PART B*/
`timescale 1ns / 1ps

module FourDigitLEDdriver(button, reset, clk, an3, an2, an1, an0, a, b, c, d, e, f, g, dp);
input clk, reset, button;
output an3, an2, an1, an0;
output a, b, c, d, e, f, g, dp;

//Set the output clks as wires:
wire clkf, clk_out, clk_outb;
reg [3:0] message [0:15];
//wire [3:0] message_w [15:0];
reg [3:0] char;

assign dp = 1'b1;

always@ (posedge clk_out or posedge reset)
begin
    if(reset) begin
        message[0] <= 4'h0;
        message[1] <= 4'h1;
        message[2] <= 4'h2;
        message[3] <= 4'h3;
        message[4] <= 4'h4;
        message[5] <= 4'h5;
        message[6] <= 4'h6;
        message[7] <= 4'h7;
        message[8] <= 4'h8;
        message[9] <= 4'h9;
        message[10] <= 4'ha;
        message[11] <= 4'hb;
        message[12] <= 4'hc;
        message[13] <= 4'hd;
        message[14] <= 4'he;
        message[15] <= 4'hf;
    end
    else begin
        message[0] <= 4'h0;
        message[1] <= 4'h1;
        message[2] <= 4'h2;
        message[3] <= 4'h3;
        message[4] <= 4'h4;
        message[5] <= 4'h5;
        message[6] <= 4'h6;
        message[7] <= 4'h7;
        message[8] <= 4'h8;
        message[9] <= 4'h9;
        message[10] <= 4'ha;
        message[11] <= 4'hb;
        message[12] <= 4'hc;
        message[13] <= 4'hd;
        message[14] <= 4'he;
        message[15] <= 4'hf;
    end
end


// MMCME2_BASE : In order to incorporate this function into the design,
//   Verilog   : the following instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (MMCME2_BASE_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // MMCME2_BASE: Base Mixed Mode Clock Manager
   //              Artix-7
   // Xilinx HDL Language Template, version 2018.3

   MMCME2_BASE #(
      .BANDWIDTH("OPTIMIZED"),   // Jitter programming (OPTIMIZED, HIGH, LOW)
      .CLKFBOUT_MULT_F(6.0),     // Multiply value for all CLKOUT (2.000-64.000).
      .CLKFBOUT_PHASE(0.0),      // Phase offset in degrees of CLKFB (-360.000-360.000).
      .CLKIN1_PERIOD(10.0),       // Input clock period in ns to ps resolution (i.e. 33.333 is 30 MHz).
      // CLKOUT0_DIVIDE - CLKOUT6_DIVIDE: Divide amount for each CLKOUT (1-128)
      .CLKOUT1_DIVIDE(120),
      .CLKOUT2_DIVIDE(1),
      .CLKOUT3_DIVIDE(1),
      .CLKOUT4_DIVIDE(1),
      .CLKOUT5_DIVIDE(1),
      .CLKOUT6_DIVIDE(1),
      .CLKOUT0_DIVIDE_F(1.0),    // Divide amount for CLKOUT0 (1.000-128.000).
      // CLKOUT0_DUTY_CYCLE - CLKOUT6_DUTY_CYCLE: Duty cycle for each CLKOUT (0.01-0.99).
      .CLKOUT0_DUTY_CYCLE(0.5),
      .CLKOUT1_DUTY_CYCLE(0.5),
      .CLKOUT2_DUTY_CYCLE(0.5),
      .CLKOUT3_DUTY_CYCLE(0.5),
      .CLKOUT4_DUTY_CYCLE(0.5),
      .CLKOUT5_DUTY_CYCLE(0.5),
      .CLKOUT6_DUTY_CYCLE(0.5),
      // CLKOUT0_PHASE - CLKOUT6_PHASE: Phase offset for each CLKOUT (-360.000-360.000).
      .CLKOUT0_PHASE(0.0),
      .CLKOUT1_PHASE(0.0),
      .CLKOUT2_PHASE(0.0),
      .CLKOUT3_PHASE(0.0),
      .CLKOUT4_PHASE(0.0),
      .CLKOUT5_PHASE(0.0),
      .CLKOUT6_PHASE(0.0),
      .CLKOUT4_CASCADE("FALSE"), // Cascade CLKOUT4 counter with CLKOUT6 (FALSE, TRUE)
      .DIVCLK_DIVIDE(1.0),         // Master division value (1-106)
      .REF_JITTER1(0.0),         // Reference input jitter in UI (0.000-0.999).
      .STARTUP_WAIT("FALSE")     // Delays DONE until MMCM is locked (FALSE, TRUE)
   )
   MMCME2_BASE_inst (
      // Clock Outputs: 1-bit (each) output: User configurable clock outputs
      .CLKOUT0(),     // 1-bit output: CLKOUT0
      .CLKOUT0B(),   // 1-bit output: Inverted CLKOUT0
      .CLKOUT1(clk_out),     // 1-bit output: CLKOUT1
      .CLKOUT1B(clk_outb),   // 1-bit output: Inverted CLKOUT1
      .CLKOUT2(),     // 1-bit output: CLKOUT2
      .CLKOUT2B(),   // 1-bit output: Inverted CLKOUT2
      .CLKOUT3(),     // 1-bit output: CLKOUT3
      .CLKOUT3B(),   // 1-bit output: Inverted CLKOUT3
      .CLKOUT4(),     // 1-bit output: CLKOUT4
      .CLKOUT5(),     // 1-bit output: CLKOUT5
      .CLKOUT6(),     // 1-bit output: CLKOUT6
      // Feedback Clocks: 1-bit (each) output: Clock feedback ports
      .CLKFBOUT(clkf),   // 1-bit output: Feedback clock
      .CLKFBOUTB(), // 1-bit output: Inverted CLKFBOUT
      // Status Ports: 1-bit (each) output: MMCM status ports
      .LOCKED(),       // 1-bit output: LOCK
      // Clock Inputs: 1-bit (each) input: Clock input
      .CLKIN1(clk),       // 1-bit input: Clock
      // Control Ports: 1-bit (each) input: MMCM control ports
      .PWRDWN(1'b0),       // 1-bit input: Power-down
      .RST(RST),             // 1-bit input: Reset
      // Feedback Clocks: 1-bit (each) input: Clock feedback ports
      .CLKFBIN(clkf)      // 1-bit input: Feedback clock
   );


integer i = 0, i0=0, i1=0, i2=0, i3=0;
reg [3:0] count;
reg en;
reg [7:0] count5;

//counter23bit counter23bit_inst(.clk(clk_out), .reset(reset), .enable(en));
always @ (posedge clk_out or posedge reset) begin  
	if (reset)  
		count5 <= 0;  
    else  
	begin
		count5 <= count5 + 1;
	end
end

always@ (posedge clk_out or posedge reset) begin  
	if(reset)
		en<=0;
	else begin
		if(count5 < 239)
			en <=1;
		else
			en <=0;
	end
end


always @ (posedge clk_out or posedge reset) begin
	if (reset)  
		char <= 0;  
    else  begin
		if(en) begin
			if((!an0)) begin
				char <= message[0+i0];
				i=i0;
				/*i0=i0+1;
				if(i0>15) 
					i0=0;*/
			end
			else if((!an1)) begin
				char <= message[1+i1];
				i=i1+1;
				/*i1=i1+1;
				if(i1>14) 
					i1=-1;*/
			end			
			else if((!an2)) begin
				char <= message[2+i2];
				i=i2+2;
				/*i2=i2+1;
				if(i2>13) 
					i2=-2;*/
			end
			else if((!an3)) begin
				char <= message[3+i3];
				i=i3+3;
				/*i3=i3+1;
				if(i3>12) 
					i3=-3;*/
			end
			else begin
				char<=message[i];
			end
		end
	   else begin
		  if((!an0)) begin
				char <= message[0+i0];
				i=i0;
				i0=i0+1;
				if(i0>15) 
					i0=0;
			end
			else if((!an1)) begin
				char <= message[1+i1];
				i=i1+1;
				i1=i1+1;
				if(i1>14) 
					i1=-1;
			end			
			else if((!an2)) begin
				char <= message[2+i2];
				i=i2+2;
				i2=i2+1;
				if(i2>13) 
					i2=-2;
			end
			else if((!an3)) begin
				char <= message[3+i3];
				i=i3+3;
				i3=i3+1;
				if(i3>12) 
					i3=-3;
			end
			else begin
				char<=message[i];
			end
	   end
    end
end


counter4bit counter4bit_inst (.clk(clk_out), .reset(reset), .an({an3, an2, an1, an0}));
LEDdecoder LEDdecoder_inst (char, {a, b, c, d, e, f, g});

endmodule